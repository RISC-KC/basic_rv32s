`ifndef STORE_VH
`define STORE_VH

`define STORE_SB 3'b000
`define STORE_SH 3'b001
`define STORE_SW 3'b010

`endif // STORE_VH