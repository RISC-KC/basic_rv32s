`ifndef RF_WD_SELECT_VH
`define RF_WD_SELECT_VH

`define RF_WD_NONE	3'b000
`define RF_WD_LOAD	3'b001
`define RF_WD_ALU	3'b010
`define RF_WD_CSR	3'b011
`define RF_WD_LUI	3'b100
`define RF_WD_JUMP	3'b101

`endif // RF_WD_SELECT_VH