`ifndef ITYPE_VH
`define ITYPE_VH

`define ITYPE_ADDI  3'b000
`define ITYPE_SLLI  3'b001
`define ITYPE_SLTI  3'b010
`define ITYPE_SLTIU 3'b011
`define ITYPE_XORI  3'b100
`define ITYPE_SRXI  3'b101
`define ITYPE_ORI   3'b110
`define ITYPE_ANDI  3'b111

`endif // ITYPE_VH