`ifndef LOAD_VH
`define LOAD_VH

`define LOAD_LB	3'b000
`define LOAD_LH	3'b001
`define LOAD_LW	3'b010
`define LOAD_LBU 3'b100
`define LOAD_LHU 3'b101

`endif // LOAD_VH