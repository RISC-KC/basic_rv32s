`ifndef TRAP_VH
`define TRAP_VH

`define TRAP_NONE		2'b00
`define TRAP_EBREAK		2'b01
`define TRAP_ECALL		2'b10
`define TRAP_MISALIGNED	2'b11

`endif // TRAP_VH