`include "modules/headers/opcode.vh"
`include "modules/headers/branch.vh"

module ALUControl (
    input [6:0] opcode,        		// opcode
	input [2:0] funct3,				// funct3
    input funct7_5,					// 5th index of funct7 (starting from 0th index)
    input imm_10,					// 10th index of imm (starting from 0th index)
	
    output reg [3:0] alu_op		// ALU operation signal
);

    always @(*) begin
        case (opcode)
			`OPCODE_RTYPE: begin
                case (funct3)
					3'b000: begin // add or sub
						alu_op = {3'b000, funct7_5};
						// add : 000 ; 0000000 
						// sub : 000 ; 0100000
					end
					3'b001: begin // sll
						alu_op = 4'b0111; // sll : 001 ; 0000000 
					end
					3'b010: begin // slt
						alu_op = 4'b0101; // slt : 010 ; 0000000
					end
					3'b011: begin // sltu
						alu_op = 4'b0110; // sltu : 011 ; 0000000
					end
					3'b100: begin // xor
						alu_op = 4'b0100; // xor : 100 ; 0000000 
					end
					3'b101: begin // srl or sra
						alu_op = {3'b100, funct7_5};
						// srl : 101 ; 0000000
						// sra : 101 ; 0100000 
					end
					3'b110: begin // or
						alu_op = 4'b0011; // or : 110 ; 0000000
					end
					3'b111: begin // and
						alu_op = 4'b0010; // and : 111 ; 0000000
					end
				endcase
            end
			`OPCODE_ITYPE: begin
				case (funct3)
					3'b000: begin
						alu_op = 4'b0000; // addi : 000 ; - 
					end
					3'b001: begin
						alu_op = 4'b0111; // slli : 001 ; imm[5:11]=0000000 
					end
					3'b010: begin
						alu_op = 4'b0101; // slti : 010 ; - 
					end
					3'b011: begin
						alu_op = 4'b0110; // sltiu : 011 ; -
					end
					3'b100: begin
						alu_op = 4'b0100; // xori : 100 ; - 
					end
					3'b101: begin
						alu_op = {3'b100, imm_10};
						// srli : 101 ; imm[5:11]=0000000 
						// srai : 101 ; imm[5:11]=0100000 
					end
					3'b110: begin
						alu_op = 4'b0011; // ori : 110 ; - 
					end
					3'b111: begin
						alu_op = 4'b0010; // andi : 111 ; -
					end
				endcase
			end
			`OPCODE_LOAD: begin
				alu_op = 4'b0000; // Every load instruction requires addition
			end
			`OPCODE_JALR: begin
				alu_op = 4'b0000; // jalr : 000 ; -
			end
			`OPCODE_STORE: begin
				alu_op = 4'b0000; // Every store instruction requires addition
			end
			`OPCODE_BRANCH: begin
				case (funct3)
					`BRANCH_BEQ: begin
						alu_op = 4'b0001; // If subtraction result is zero, equal
					end
					`BRANCH_BNE: begin
						alu_op = 4'b0001; // If subtraction result is not zero, not equal
					end
					`BRANCH_BLT: begin
						alu_op = 4'b0101; // If SLT result is not zero, less
					end
					`BRANCH_BGE: begin
						alu_op = 4'b0101; // If SLT result is zero, greater or equal
					end
					`BRANCH_BLTU: begin
						alu_op = 4'b0110; // If SLTU result is not zero, less (unsigned)
					end
					`BRANCH_BGEU: begin
						alu_op = 4'b0110; // If SLTU result is zero, greater or equal (unsigned)
					end
				endcase
			end
			`OPCODE_ENVIRONMENT: begin
				case (funct3)
					3'b001: begin // csrrw : 001 ; -
						alu_op = 4'b1111;
					end
					3'b010: begin // csrrs : 010 ; -
						alu_op = 4'b0011;
					end
					3'b011: begin // csrrc : 011 ; -
						alu_op = 4'b1010;
					end
					3'b101: begin // csrrwi : 101 ; -
						alu_op = 4'b1111;
					end
					3'b110: begin // csrrsi : 110 ; -
						alu_op = 4'b0011;
					end
					3'b111: begin // csrrci : 111 ; -
						alu_op = 4'b1010;
					end
					default: begin
						alu_op = 4'b1111;
					end
				endcase
			end
			default: begin
				alu_op = 4'b1111;
			end
        endcase
    end

endmodule
